module network

pub struct RPC {
pub:
	payload []u8
}
