module core

type Timestamp = u64
