module network

pub interface INetworkEndpoint {
}
